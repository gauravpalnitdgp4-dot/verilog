// -----------------------------------------------------------------------------
// Module: odd_div
// Description:
//   Parameterizable clock divider that divides the input clock (clk) by an odd or
//   even value specified by div_val. Generates clkout with ~50% duty cycle for
//   both odd and even division values.
//
// Ports:
//   input  logic resetn   - Active-low reset. Resets all internal registers.
//   input  logic [7:0] div_val - Division value (odd/even supported).
//   input  logic clk      - Input clock to be divided.
//   output logic clkout   - Output divided clock.
//
// Internal Signals:
//   logic [7:0] cnt       - Counts clock cycles up to div_val - 1.
//   logic toggle1, toggle2- Toggles for generating clkout with correct duty cycle.
//   logic [6:0] half_div  - Half of div_val (integer division).
//   logic odd_even        - 1 if div_val is odd, 0 if even.
//   logic [7:0] div_val_lat - Latched division value for stable operation.
//
// Functionality:
//   - On reset, all signals are initialized.
//   - div_val is latched at the start of each division cycle.
//   - For odd div_val: toggle1 toggles every div_val cycles, toggle2 toggles at midpoint.
//   - For even div_val: toggle1 toggles every div_val/2 cycles.
//   - clkout is generated by combining toggle1 and toggle2 for odd division, or just toggle1 for even division.
//
// Output Logic:
//   clkout = (odd_even) ? (toggle1 ^ toggle2) : toggle1;
// -----------------------------------------------------------------------------

module odd_div (
    input logic resetn,
    input logic [7:0] div_val,
    input logic clk,
    output logic clkout
);
    logic [7:0] cnt;
    logic toggle1;
    logic toggle2;
    logic [6:0] half_div;
    logic odd_even;
    logic [7:0] div_val_lat;
    assign half_div = (cnt == 0)? div_val[7:1]: div_val_lat[7:1]; // Integer division by 2
    assign odd_even = (cnt == 0)? div_val[0]: div_val_lat[0]; // 1 if odd, 0 if even
    // For odd div_val, toggle1 toggles every div_val cycles
    // For even div_val, toggle1 toggles every div_val/2 cycles
    always_ff @(posedge clk or negedge resetn) begin
        if (!resetn) begin
            div_val_lat <= 0;
        end else if (cnt == 0) begin
            div_val_lat <= div_val;
        end
    end
    always_ff @(posedge clk or negedge resetn) begin
        if (!resetn) begin
            cnt <= 0;
            toggle1 <= 1;
            toggle2 <= 1;
        end else begin 
            if (cnt == 0 & odd_even == 1'b1) begin
                toggle1 <= ~toggle1;
            end
            else if (((cnt == 0)|cnt == (half_div))  & odd_even == 1'b0) begin
                toggle1 <= ~toggle1;
            end
            cnt <= (cnt == div_val_lat - 1) ? 0 : cnt + 1;
        end
    end
    always_ff @(negedge clk or negedge resetn) begin
        if (!resetn) begin
            toggle2 <= 1;
        end else begin 
            if (cnt == (half_div + 1)) begin
                toggle2 <= ~toggle2;
            end
        end
    end
assign clkout = (odd_even) ? (toggle1 ^ toggle2) : toggle1;
endmodule

